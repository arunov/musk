package CACHE;

typedef enum { READ, WRITE } cmd_t;

endpackage
