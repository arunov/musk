package CACHE;

typedef enum {IDLE, READ, WRITE, FLUSH} cache_cmd_t;

endpackage
