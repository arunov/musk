
module MPipeline(
);

endmodule
