package DECODER;

`include "DecoderTypes.sv"
`include "OpcodeMap.sv"
`include "OperandDecoder.sv"
`include "Decoder.sv"

endpackage
