
import DecoderTypes::*;

module APipeline(
	input logic reset,
	input logic clk,
);

endmodule
