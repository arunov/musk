package DECODER;

`include "DecoderTypes.sv"
`include "OpcodeMap.sv"
`include "OperandDecoder.sv"
`include "MainDecoder.sv"

endpackage
