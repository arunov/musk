package MicroOp;

import DecoderTypes::*;


endpackage
