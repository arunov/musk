package InstructionPrinter;

import DecoderTypes::*;
import RegMap::*;

endpackage
